tyler is a gooner
