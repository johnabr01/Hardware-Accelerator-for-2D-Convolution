`define INWVAL 12
`define RVAL 9
`define CVAL 8
`define MAXKVAL 5
`define TVPR 1
`define TRPR 1
