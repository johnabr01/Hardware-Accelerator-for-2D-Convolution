blahahah